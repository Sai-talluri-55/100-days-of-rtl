`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.12.2023 19:05:30
// Design Name: 
// Module Name: johnsoncounter_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module johnsoncounter_tb(

    );
    reg clk,rst;
wire [3:0]q;
johnson_counter dut(clk,rst,q);
initial clk=0;
always #5 clk=~clk;
initial 
begin
rst=1;
#20 rst=0;
#100 $finish;
end
endmodule
